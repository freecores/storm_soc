-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 15.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
				MEM_SIZE      : natural := 1024;  -- memory cells
				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
		000000 => x"EA000006",
		000001 => x"EAFFFFFE",
		000002 => x"EAFFFFFE",
		000003 => x"EAFFFFFE",
		000004 => x"EAFFFFFE",
		000005 => x"E1A00000",
		000006 => x"EAFFFFFE",
		000007 => x"EAFFFFFE",
		000008 => x"E59F0034",
		000009 => x"E10F1000",
		000010 => x"E3C1107F",
		000011 => x"E38110DF",
		000012 => x"E129F001",
		000013 => x"E1A0D000",
		000014 => x"E3A00000",
		000015 => x"E1A01000",
		000016 => x"E1A02000",
		000017 => x"E1A0B000",
		000018 => x"E1A07000",
		000019 => x"E59FA00C",
		000020 => x"E1A0E00F",
		000021 => x"E1A0F00A",
		000022 => x"EAFFFFFE",
		000023 => x"00008000",
		000024 => x"FFF00700",
		000025 => x"E3E03A0F",
		000026 => x"E5131FFB",
		000027 => x"E20020FF",
		000028 => x"E3A00001",
		000029 => x"E0010210",
		000030 => x"E1A0F00E",
		000031 => x"E3E03A0F",
		000032 => x"E5130FFB",
		000033 => x"E1A0F00E",
		000034 => x"E3E01A0F",
		000035 => x"E5113FFF",
		000036 => x"E20000FF",
		000037 => x"E3A02001",
		000038 => x"E1833012",
		000039 => x"E5013FFF",
		000040 => x"E1A0F00E",
		000041 => x"E20000FF",
		000042 => x"E3A02001",
		000043 => x"E1A02012",
		000044 => x"E3E01A0F",
		000045 => x"E5113FFF",
		000046 => x"E1E02002",
		000047 => x"E0033002",
		000048 => x"E5013FFF",
		000049 => x"E1A0F00E",
		000050 => x"E3E01A0F",
		000051 => x"E5113FFF",
		000052 => x"E20000FF",
		000053 => x"E3A02001",
		000054 => x"E0233012",
		000055 => x"E5013FFF",
		000056 => x"E1A0F00E",
		000057 => x"E3E03A0F",
		000058 => x"E5030FFF",
		000059 => x"E1A0F00E",
		000060 => x"E20000FF",
		000061 => x"E3500007",
		000062 => x"E92D4010",
		000063 => x"E3A0C000",
		000064 => x"E3E0E0FF",
		000065 => x"E20110FF",
		000066 => x"8A000011",
		000067 => x"E2403004",
		000068 => x"E20330FF",
		000069 => x"E3500003",
		000070 => x"E1A0E183",
		000071 => x"E3E04A0F",
		000072 => x"E1A0C180",
		000073 => x"9A000007",
		000074 => x"E3A030FF",
		000075 => x"E1A03E13",
		000076 => x"E5142F8B",
		000077 => x"E1E03003",
		000078 => x"E0022003",
		000079 => x"E1822E11",
		000080 => x"E5042F8B",
		000081 => x"E8BD8010",
		000082 => x"E3A030FF",
		000083 => x"E1A03C13",
		000084 => x"E1E0E003",
		000085 => x"E3E02A0F",
		000086 => x"E5123F8F",
		000087 => x"E003300E",
		000088 => x"E1833C11",
		000089 => x"E5023F8F",
		000090 => x"E8BD8010",
		000091 => x"E20000FF",
		000092 => x"E3500007",
		000093 => x"E3A02000",
		000094 => x"8A00000A",
		000095 => x"E2403004",
		000096 => x"E3500003",
		000097 => x"E20320FF",
		000098 => x"9A000005",
		000099 => x"E3E03A0F",
		000100 => x"E5130F8B",
		000101 => x"E1A02182",
		000102 => x"E1A00230",
		000103 => x"E20000FF",
		000104 => x"E1A0F00E",
		000105 => x"E1A02180",
		000106 => x"E3E03A0F",
		000107 => x"E5130F8F",
		000108 => x"E1A00230",
		000109 => x"E20000FF",
		000110 => x"E1A0F00E",
		000111 => x"E3E02A0F",
		000112 => x"E5123FE3",
		000113 => x"E3130002",
		000114 => x"E3E00000",
		000115 => x"15120FE7",
		000116 => x"E1A0F00E",
		000117 => x"E3E02A0F",
		000118 => x"E5123FE3",
		000119 => x"E3130001",
		000120 => x"0AFFFFFC",
		000121 => x"E20030FF",
		000122 => x"E5023FE7",
		000123 => x"E1A0F00E",
		000124 => x"E20000FF",
		000125 => x"E3500001",
		000126 => x"E3812B01",
		000127 => x"03E03A0F",
		000128 => x"E3811B09",
		000129 => x"13E03A0F",
		000130 => x"05031FCF",
		000131 => x"15032FCF",
		000132 => x"E1A0F00E",
		000133 => x"E3E03A0F",
		000134 => x"E5030FCB",
		000135 => x"E1A0F00E",
		000136 => x"E3E02A0F",
		000137 => x"E5123FCF",
		000138 => x"E3130C01",
		000139 => x"1AFFFFFC",
		000140 => x"E5020FBF",
		000141 => x"E5123FCF",
		000142 => x"E3833C01",
		000143 => x"E5023FCF",
		000144 => x"E3E02A0F",
		000145 => x"E5123FCF",
		000146 => x"E3130C01",
		000147 => x"1AFFFFFC",
		000148 => x"E5120FBF",
		000149 => x"E1A0F00E",
		000150 => x"E3E01A0F",
		000151 => x"E5113FC7",
		000152 => x"E20000FF",
		000153 => x"E3A02001",
		000154 => x"E1833012",
		000155 => x"E5013FC7",
		000156 => x"E1A0F00E",
		000157 => x"E20000FF",
		000158 => x"E3A02001",
		000159 => x"E1A02012",
		000160 => x"E3E01A0F",
		000161 => x"E5113FC7",
		000162 => x"E1E02002",
		000163 => x"E0033002",
		000164 => x"E5013FC7",
		000165 => x"E1A0F00E",
		000166 => x"E3E02A0F",
		000167 => x"E5123F97",
		000168 => x"E1A01420",
		000169 => x"E3C33080",
		000170 => x"E5023F97",
		000171 => x"E5020F9F",
		000172 => x"E5021F9B",
		000173 => x"E5123F97",
		000174 => x"E3833080",
		000175 => x"E5023F97",
		000176 => x"E1A0F00E",
		000177 => x"E92D4030",
		000178 => x"E3A0C090",
		000179 => x"E20140FE",
		000180 => x"E3E0EA0F",
		000181 => x"E5DD500F",
		000182 => x"E20000FF",
		000183 => x"E50E4F93",
		000184 => x"E20110FF",
		000185 => x"E50ECFAF",
		000186 => x"E1A04002",
		000187 => x"E203C0FF",
		000188 => x"E51E3FAF",
		000189 => x"E3130002",
		000190 => x"1AFFFFFC",
		000191 => x"E51E3FAF",
		000192 => x"E3130080",
		000193 => x"13E00000",
		000194 => x"18BD8030",
		000195 => x"E35C0000",
		000196 => x"0A000012",
		000197 => x"E24C3001",
		000198 => x"E203C0FF",
		000199 => x"E35C0001",
		000200 => x"01A02424",
		000201 => x"03E03A0F",
		000202 => x"13E03A0F",
		000203 => x"05032F93",
		000204 => x"15034F93",
		000205 => x"E3E02A0F",
		000206 => x"E3A03010",
		000207 => x"E5023FAF",
		000208 => x"E5123FAF",
		000209 => x"E3130002",
		000210 => x"1AFFFFFC",
		000211 => x"E5123FAF",
		000212 => x"E3130080",
		000213 => x"0AFFFFEC",
		000214 => x"E3E00001",
		000215 => x"E8BD8030",
		000216 => x"E3500077",
		000217 => x"1A00000C",
		000218 => x"E3E03A0F",
		000219 => x"E3A02050",
		000220 => x"E5035F93",
		000221 => x"E5032FAF",
		000222 => x"E1A02003",
		000223 => x"E5123FAF",
		000224 => x"E3130002",
		000225 => x"1AFFFFFC",
		000226 => x"E5123FAF",
		000227 => x"E2130080",
		000228 => x"08BD8030",
		000229 => x"E3E00002",
		000230 => x"E8BD8030",
		000231 => x"E3500072",
		000232 => x"13E00003",
		000233 => x"18BD8030",
		000234 => x"E3813001",
		000235 => x"E3E02A0F",
		000236 => x"E3A01090",
		000237 => x"E5023F93",
		000238 => x"E5021FAF",
		000239 => x"E5123FAF",
		000240 => x"E3130002",
		000241 => x"1AFFFFFC",
		000242 => x"E5123FAF",
		000243 => x"E3130080",
		000244 => x"1AFFFFEF",
		000245 => x"E3A03068",
		000246 => x"E5023FAF",
		000247 => x"E3E00A0F",
		000248 => x"E5103FAF",
		000249 => x"E3130002",
		000250 => x"1AFFFFFC",
		000251 => x"E5100F93",
		000252 => x"E8BD8030",
		000253 => x"E20000FF",
		000254 => x"E350000D",
		000255 => x"979FF100",
		000256 => x"EA000015",
		000257 => x"FFF0043C",
		000258 => x"FFF00484",
		000259 => x"FFF0047C",
		000260 => x"FFF0045C",
		000261 => x"FFF0045C",
		000262 => x"FFF0045C",
		000263 => x"FFF00474",
		000264 => x"FFF0045C",
		000265 => x"FFF0046C",
		000266 => x"FFF00464",
		000267 => x"FFF0045C",
		000268 => x"FFF00454",
		000269 => x"FFF0044C",
		000270 => x"FFF00444",
		000271 => x"EE100F10",
		000272 => x"E1A0F00E",
		000273 => x"EE1D0F1D",
		000274 => x"E1A0F00E",
		000275 => x"EE1C0F1C",
		000276 => x"E1A0F00E",
		000277 => x"EE1B0F1B",
		000278 => x"E1A0F00E",
		000279 => x"E3A00000",
		000280 => x"E1A0F00E",
		000281 => x"EE190F19",
		000282 => x"E1A0F00E",
		000283 => x"EE180F18",
		000284 => x"E1A0F00E",
		000285 => x"EE160F16",
		000286 => x"E1A0F00E",
		000287 => x"EE120F12",
		000288 => x"E1A0F00E",
		000289 => x"EE110F11",
		000290 => x"E1A0F00E",
		000291 => x"E20110FF",
		000292 => x"E2411006",
		000293 => x"E3510007",
		000294 => x"979FF101",
		000295 => x"EA000008",
		000296 => x"FFF004C8",
		000297 => x"FFF004C4",
		000298 => x"FFF004C4",
		000299 => x"FFF004C4",
		000300 => x"FFF004C4",
		000301 => x"FFF004D0",
		000302 => x"FFF004D8",
		000303 => x"FFF004C0",
		000304 => x"EE0D0F1D",
		000305 => x"E1A0F00E",
		000306 => x"EE060F16",
		000307 => x"E1A0F00E",
		000308 => x"EE0B0F1B",
		000309 => x"E1A0F00E",
		000310 => x"EE0C0F1C",
		000311 => x"E1A0F00E",
		000312 => x"E10F0000",
		000313 => x"E1A0F00E",
		000314 => x"E129F000",
		000315 => x"E1A0F00E",
		000316 => x"E52DE004",
		000317 => x"EBFFFFF9",
		000318 => x"E3C00080",
		000319 => x"E49DE004",
		000320 => x"EAFFFFF8",
		000321 => x"E52DE004",
		000322 => x"EBFFFFF4",
		000323 => x"E3800080",
		000324 => x"E49DE004",
		000325 => x"EAFFFFF3",
		000326 => x"E92D4010",
		000327 => x"E1A04000",
		000328 => x"E5D00000",
		000329 => x"E3500000",
		000330 => x"1A000003",
		000331 => x"EA000005",
		000332 => x"E5F40001",
		000333 => x"E3500000",
		000334 => x"0A000002",
		000335 => x"EBFFFF24",
		000336 => x"E3500000",
		000337 => x"CAFFFFF9",
		000338 => x"E1A00004",
		000339 => x"E8BD8010",
		000340 => x"E92D4070",
		000341 => x"E2514000",
		000342 => x"E1A05000",
		000343 => x"E20260FF",
		000344 => x"D8BD8070",
		000345 => x"EBFFFF14",
		000346 => x"E3700001",
		000347 => x"E20030FF",
		000348 => x"0A000005",
		000349 => x"E3560001",
		000350 => x"E5C53000",
		000351 => x"E1A00003",
		000352 => x"E2855001",
		000353 => x"0A000003",
		000354 => x"E2444001",
		000355 => x"E3540000",
		000356 => x"CAFFFFF3",
		000357 => x"E8BD8070",
		000358 => x"EBFFFF0D",
		000359 => x"EAFFFFF9",
		000360 => x"E92D4030",
		000361 => x"E2514000",
		000362 => x"E1A05000",
		000363 => x"D8BD8030",
		000364 => x"E4D50001",
		000365 => x"EBFFFF06",
		000366 => x"E2544001",
		000367 => x"1AFFFFFB",
		000368 => x"E8BD8030",
		000369 => x"E92D4010",
		000370 => x"E20240FF",
		000371 => x"E3540008",
		000372 => x"83A04008",
		000373 => x"8A000001",
		000374 => x"E3540000",
		000375 => x"03A04001",
		000376 => x"E1A02001",
		000377 => x"E1A0E004",
		000378 => x"E1A0310E",
		000379 => x"E35E0001",
		000380 => x"E2433004",
		000381 => x"E1A0C000",
		000382 => x"81A0C330",
		000383 => x"E24E3001",
		000384 => x"E20CC00F",
		000385 => x"E203E0FF",
		000386 => x"E35C0009",
		000387 => x"E28C3030",
		000388 => x"828C3037",
		000389 => x"E35E0000",
		000390 => x"E4C23001",
		000391 => x"1AFFFFF1",
		000392 => x"E2443001",
		000393 => x"E20330FF",
		000394 => x"E0813003",
		000395 => x"E5C3E001",
		000396 => x"E8BD8010",
		000397 => x"E20110FF",
		000398 => x"E3510008",
		000399 => x"E92D4010",
		000400 => x"E1A04000",
		000401 => x"8A000016",
		000402 => x"E3510000",
		000403 => x"0A000014",
		000404 => x"E3A00000",
		000405 => x"EA000006",
		000406 => x"E2413001",
		000407 => x"E20310FF",
		000408 => x"E202200F",
		000409 => x"E1A03101",
		000410 => x"E3510000",
		000411 => x"E1800312",
		000412 => x"08BD8010",
		000413 => x"E4D43001",
		000414 => x"E2432030",
		000415 => x"E3520009",
		000416 => x"E243C041",
		000417 => x"9AFFFFF3",
		000418 => x"E35C0005",
		000419 => x"E243E061",
		000420 => x"E2432037",
		000421 => x"9AFFFFEF",
		000422 => x"E35E0005",
		000423 => x"E2432057",
		000424 => x"9AFFFFEC",
		000425 => x"E3A00000",
		000426 => x"E8BD8010",
		000427 => x"E1A03000",
		000428 => x"E5D00001",
		000429 => x"E283C001",
		000430 => x"E5D32000",
		000431 => x"E5DC1002",
		000432 => x"E1A00800",
		000433 => x"E1800C02",
		000434 => x"E5DC3001",
		000435 => x"E1800001",
		000436 => x"E1800403",
		000437 => x"E1A0F00E",
		000438 => x"E0603280",
		000439 => x"E0800103",
		000440 => x"E0800100",
		000441 => x"E1A00200",
		000442 => x"E3500000",
		000443 => x"D1A0F00E",
		000444 => x"E1A00000",
		000445 => x"E2500001",
		000446 => x"1AFFFFFC",
		000447 => x"E1A0F00E",
		000448 => x"E92D45F0",
		000449 => x"E3A00000",
		000450 => x"E24DD00C",
		000451 => x"EBFFFE74",
		000452 => x"E3A0100D",
		000453 => x"E3A000C3",
		000454 => x"EBFFFF5B",
		000455 => x"E3A00063",
		000456 => x"EBFFFEDC",
		000457 => x"E3A00006",
		000458 => x"EBFFFF31",
		000459 => x"E3A01006",
		000460 => x"E3800008",
		000461 => x"EBFFFF54",
		000462 => x"E3A0000D",
		000463 => x"EBFFFF2C",
		000464 => x"E1A000A0",
		000465 => x"E1E00000",
		000466 => x"E200000F",
		000467 => x"E3500001",
		000468 => x"028DA007",
		000469 => x"0A00001B",
		000470 => x"E3500002",
		000471 => x"02800001",
		000472 => x"028DA007",
		000473 => x"0A000017",
		000474 => x"E59F0934",
		000475 => x"EBFFFF69",
		000476 => x"E59F0930",
		000477 => x"EBFFFF67",
		000478 => x"E59F092C",
		000479 => x"EBFFFF65",
		000480 => x"E59F0928",
		000481 => x"EBFFFF63",
		000482 => x"E59F0924",
		000483 => x"EBFFFF61",
		000484 => x"E59F0920",
		000485 => x"EBFFFF5F",
		000486 => x"E59F091C",
		000487 => x"EBFFFF5D",
		000488 => x"E59F0918",
		000489 => x"EBFFFF5B",
		000490 => x"E59F0914",
		000491 => x"EBFFFF59",
		000492 => x"E59F0910",
		000493 => x"EBFFFF57",
		000494 => x"E59F090C",
		000495 => x"EBFFFF55",
		000496 => x"E28DA007",
		000497 => x"EBFFFE7C",
		000498 => x"E2803001",
		000499 => x"E3530073",
		000500 => x"979FF103",
		000501 => x"EA0001AF",
		000502 => x"FFF009E8",
		000503 => x"FFF00E98",
		000504 => x"FFF00E98",
		000505 => x"FFF00E98",
		000506 => x"FFF00E98",
		000507 => x"FFF00E98",
		000508 => x"FFF00E98",
		000509 => x"FFF00E98",
		000510 => x"FFF00E98",
		000511 => x"FFF00E98",
		000512 => x"FFF00E98",
		000513 => x"FFF00E98",
		000514 => x"FFF00E98",
		000515 => x"FFF00E98",
		000516 => x"FFF00E98",
		000517 => x"FFF00E98",
		000518 => x"FFF00E98",
		000519 => x"FFF00E98",
		000520 => x"FFF00E98",
		000521 => x"FFF00E98",
		000522 => x"FFF00E98",
		000523 => x"FFF00E98",
		000524 => x"FFF00E98",
		000525 => x"FFF00E98",
		000526 => x"FFF00E98",
		000527 => x"FFF00E98",
		000528 => x"FFF00E98",
		000529 => x"FFF00E98",
		000530 => x"FFF00E98",
		000531 => x"FFF00E98",
		000532 => x"FFF00E98",
		000533 => x"FFF00E98",
		000534 => x"FFF00E98",
		000535 => x"FFF00E98",
		000536 => x"FFF00E98",
		000537 => x"FFF00E98",
		000538 => x"FFF00E98",
		000539 => x"FFF00E98",
		000540 => x"FFF00E98",
		000541 => x"FFF00E98",
		000542 => x"FFF00E98",
		000543 => x"FFF00E98",
		000544 => x"FFF00E98",
		000545 => x"FFF00E98",
		000546 => x"FFF00E98",
		000547 => x"FFF00E98",
		000548 => x"FFF00E98",
		000549 => x"FFF00E98",
		000550 => x"FFF00E98",
		000551 => x"FFF00A28",
		000552 => x"FFF00A34",
		000553 => x"FFF00AEC",
		000554 => x"FFF00B60",
		000555 => x"FFF00D38",
		000556 => x"FFF00D78",
		000557 => x"FFF00E98",
		000558 => x"FFF00E98",
		000559 => x"FFF00E98",
		000560 => x"FFF00E98",
		000561 => x"FFF00E98",
		000562 => x"FFF00E98",
		000563 => x"FFF00E98",
		000564 => x"FFF00E98",
		000565 => x"FFF00E98",
		000566 => x"FFF00E98",
		000567 => x"FFF00E98",
		000568 => x"FFF00E98",
		000569 => x"FFF00E98",
		000570 => x"FFF00E98",
		000571 => x"FFF00E98",
		000572 => x"FFF00E98",
		000573 => x"FFF00E98",
		000574 => x"FFF00E98",
		000575 => x"FFF00E98",
		000576 => x"FFF00E98",
		000577 => x"FFF00E98",
		000578 => x"FFF00E98",
		000579 => x"FFF00E98",
		000580 => x"FFF00E98",
		000581 => x"FFF00E98",
		000582 => x"FFF00E98",
		000583 => x"FFF00E98",
		000584 => x"FFF00E98",
		000585 => x"FFF00E98",
		000586 => x"FFF00E98",
		000587 => x"FFF00E98",
		000588 => x"FFF00E98",
		000589 => x"FFF00E98",
		000590 => x"FFF00E98",
		000591 => x"FFF00E98",
		000592 => x"FFF00E98",
		000593 => x"FFF00E98",
		000594 => x"FFF00E98",
		000595 => x"FFF00E98",
		000596 => x"FFF00E98",
		000597 => x"FFF00E98",
		000598 => x"FFF00E98",
		000599 => x"FFF00E98",
		000600 => x"FFF00EC0",
		000601 => x"FFF00E98",
		000602 => x"FFF00E98",
		000603 => x"FFF00E98",
		000604 => x"FFF00E98",
		000605 => x"FFF00EE4",
		000606 => x"FFF00E98",
		000607 => x"FFF00DB8",
		000608 => x"FFF00E64",
		000609 => x"FFF00E98",
		000610 => x"FFF00E98",
		000611 => x"FFF00E98",
		000612 => x"FFF00E98",
		000613 => x"FFF00E98",
		000614 => x"FFF00E98",
		000615 => x"FFF00E98",
		000616 => x"FFF00E98",
		000617 => x"FFF00EAC",
		000618 => x"E59F0720",
		000619 => x"EBFFFED9",
		000620 => x"E1A0000A",
		000621 => x"E3A01004",
		000622 => x"E3A02000",
		000623 => x"EBFFFEE3",
		000624 => x"E5DD3007",
		000625 => x"E3530053",
		000626 => x"1A000002",
		000627 => x"E5DD2008",
		000628 => x"E352004D",
		000629 => x"0A000169",
		000630 => x"E59F06F4",
		000631 => x"EBFFFECD",
		000632 => x"E59F06F0",
		000633 => x"EBFFFECB",
		000634 => x"E3A0000D",
		000635 => x"EBFFFE80",
		000636 => x"E3100001",
		000637 => x"1AFFFF72",
		000638 => x"E59F06DC",
		000639 => x"EBFFFEC5",
		000640 => x"E3A0100D",
		000641 => x"E3A00000",
		000642 => x"EBFFFE9F",
		000643 => x"E3A00006",
		000644 => x"EBFFFE77",
		000645 => x"E3A01006",
		000646 => x"E3C00008",
		000647 => x"EBFFFE9A",
		000648 => x"E3A0F000",
		000649 => x"EAFFFFFE",
		000650 => x"E3A00030",
		000651 => x"EBFFFDE8",
		000652 => x"EAFFFFF0",
		000653 => x"E3A00031",
		000654 => x"EBFFFDE5",
		000655 => x"E59F069C",
		000656 => x"EBFFFEB4",
		000657 => x"E1A0000A",
		000658 => x"E3A01004",
		000659 => x"E3A02000",
		000660 => x"EBFFFEBE",
		000661 => x"E5DD3007",
		000662 => x"E3530053",
		000663 => x"1A000002",
		000664 => x"E5DD3008",
		000665 => x"E353004D",
		000666 => x"0A000002",
		000667 => x"E59F0670",
		000668 => x"EBFFFEA8",
		000669 => x"EAFFFFDB",
		000670 => x"E5DD3009",
		000671 => x"E3530042",
		000672 => x"1AFFFFF9",
		000673 => x"E5DD300A",
		000674 => x"E3530052",
		000675 => x"1AFFFFF6",
		000676 => x"E3A01004",
		000677 => x"E3A02000",
		000678 => x"E1A0000A",
		000679 => x"EBFFFEAB",
		000680 => x"E1A0000A",
		000681 => x"EBFFFF00",
		000682 => x"E3A03C7F",
		000683 => x"E28330F8",
		000684 => x"E1500003",
		000685 => x"8A00009C",
		000686 => x"E2905004",
		000687 => x"0AFFFFCD",
		000688 => x"E3A04000",
		000689 => x"E3A01004",
		000690 => x"E3A02000",
		000691 => x"E1A0000A",
		000692 => x"EBFFFE9E",
		000693 => x"E1A0000A",
		000694 => x"EBFFFEF3",
		000695 => x"E4840004",
		000696 => x"E1550004",
		000697 => x"1AFFFFF6",
		000698 => x"EAFFFFC2",
		000699 => x"E3A00032",
		000700 => x"EBFFFDB7",
		000701 => x"E59F05EC",
		000702 => x"EBFFFE86",
		000703 => x"EBFFFDAE",
		000704 => x"E3700001",
		000705 => x"0AFFFFFC",
		000706 => x"EBFFFDAB",
		000707 => x"E3700001",
		000708 => x"1AFFFFFC",
		000709 => x"E3A05000",
		000710 => x"E5954000",
		000711 => x"E1A00C24",
		000712 => x"EBFFFDAB",
		000713 => x"E1A00824",
		000714 => x"EBFFFDA9",
		000715 => x"E1A00424",
		000716 => x"EBFFFDA7",
		000717 => x"E1A00004",
		000718 => x"EBFFFDA5",
		000719 => x"EBFFFD9E",
		000720 => x"E3700001",
		000721 => x"E2855004",
		000722 => x"1A000001",
		000723 => x"E3550902",
		000724 => x"1AFFFFF0",
		000725 => x"E59F0590",
		000726 => x"EBFFFE6E",
		000727 => x"EAFFFFA1",
		000728 => x"E3A04000",
		000729 => x"E59F0584",
		000730 => x"EBFFFE6A",
		000731 => x"E1A01006",
		000732 => x"E1A02004",
		000733 => x"E3A03002",
		000734 => x"E3A00072",
		000735 => x"E58D4000",
		000736 => x"EBFFFDCF",
		000737 => x"E1A01006",
		000738 => x"E5CD0007",
		000739 => x"E3A02001",
		000740 => x"E3A03002",
		000741 => x"E3A00072",
		000742 => x"E58D4000",
		000743 => x"EBFFFDC8",
		000744 => x"E3A02002",
		000745 => x"E1A03002",
		000746 => x"E5CD0008",
		000747 => x"E1A01006",
		000748 => x"E3A00072",
		000749 => x"E58D4000",
		000750 => x"EBFFFDC1",
		000751 => x"E3A03002",
		000752 => x"E5CD0009",
		000753 => x"E1A01006",
		000754 => x"E3A00072",
		000755 => x"E3A02003",
		000756 => x"E58D4000",
		000757 => x"EBFFFDBA",
		000758 => x"E5DD3007",
		000759 => x"E20000FF",
		000760 => x"E3530053",
		000761 => x"E5CD000A",
		000762 => x"1A000002",
		000763 => x"E5DD3008",
		000764 => x"E353004D",
		000765 => x"0A000002",
		000766 => x"E59F04F4",
		000767 => x"EBFFFE45",
		000768 => x"EAFFFF78",
		000769 => x"E5DD3009",
		000770 => x"E3530042",
		000771 => x"1AFFFFF9",
		000772 => x"E3500052",
		000773 => x"1AFFFFF7",
		000774 => x"E1A01006",
		000775 => x"E3A02004",
		000776 => x"E2433040",
		000777 => x"E2800020",
		000778 => x"E58D4000",
		000779 => x"EBFFFDA4",
		000780 => x"E1A01006",
		000781 => x"E5CD0007",
		000782 => x"E3A02005",
		000783 => x"E3A03002",
		000784 => x"E3A00072",
		000785 => x"E58D4000",
		000786 => x"EBFFFD9D",
		000787 => x"E1A01006",
		000788 => x"E5CD0008",
		000789 => x"E3A02006",
		000790 => x"E3A03002",
		000791 => x"E3A00072",
		000792 => x"E58D4000",
		000793 => x"EBFFFD96",
		000794 => x"E1A01006",
		000795 => x"E5CD0009",
		000796 => x"E3A02007",
		000797 => x"E3A03002",
		000798 => x"E3A00072",
		000799 => x"E58D4000",
		000800 => x"EBFFFD8F",
		000801 => x"E5CD000A",
		000802 => x"E1A0000A",
		000803 => x"EBFFFE86",
		000804 => x"E2907004",
		000805 => x"0A000021",
		000806 => x"E1A05004",
		000807 => x"E2842008",
		000808 => x"E1A01006",
		000809 => x"E3A03002",
		000810 => x"E3A00072",
		000811 => x"E58D5000",
		000812 => x"EBFFFD83",
		000813 => x"E2842009",
		000814 => x"E5CD0007",
		000815 => x"E1A01006",
		000816 => x"E3A03002",
		000817 => x"E3A00072",
		000818 => x"E58D5000",
		000819 => x"EBFFFD7C",
		000820 => x"E284200A",
		000821 => x"E5CD0008",
		000822 => x"E1A01006",
		000823 => x"E3A03002",
		000824 => x"E3A00072",
		000825 => x"E58D5000",
		000826 => x"EBFFFD75",
		000827 => x"E284200B",
		000828 => x"E5CD0009",
		000829 => x"E1A01006",
		000830 => x"E3A03002",
		000831 => x"E3A00072",
		000832 => x"E58D5000",
		000833 => x"EBFFFD6E",
		000834 => x"E5CD000A",
		000835 => x"E1A0000A",
		000836 => x"EBFFFE65",
		000837 => x"E4840004",
		000838 => x"E1540007",
		000839 => x"1AFFFFDE",
		000840 => x"E59F03D0",
		000841 => x"EBFFFDFB",
		000842 => x"EAFFFF32",
		000843 => x"E59F03C8",
		000844 => x"EBFFFDF8",
		000845 => x"EAFFFF2B",
		000846 => x"E3A00034",
		000847 => x"EBFFFD24",
		000848 => x"E59F03B8",
		000849 => x"EBFFFDF3",
		000850 => x"E1A0000A",
		000851 => x"E3A01002",
		000852 => x"E3A02001",
		000853 => x"EBFFFDFD",
		000854 => x"E1A0000A",
		000855 => x"E3A01002",
		000856 => x"EBFFFE33",
		000857 => x"E21060FF",
		000858 => x"1AFFFF0E",
		000859 => x"E59F0390",
		000860 => x"EBFFFDE8",
		000861 => x"EAFFFF1B",
		000862 => x"E3A00035",
		000863 => x"EBFFFD14",
		000864 => x"E59F0380",
		000865 => x"EBFFFDE3",
		000866 => x"E1A0000A",
		000867 => x"E3A01002",
		000868 => x"E3A02001",
		000869 => x"EBFFFDED",
		000870 => x"E1A0000A",
		000871 => x"E3A01002",
		000872 => x"EBFFFE23",
		000873 => x"E21060FF",
		000874 => x"1A000054",
		000875 => x"E59F0358",
		000876 => x"EBFFFDD8",
		000877 => x"EAFFFF0B",
		000878 => x"E3A00068",
		000879 => x"EBFFFD04",
		000880 => x"E59F0348",
		000881 => x"EBFFFDD3",
		000882 => x"E59F0344",
		000883 => x"EBFFFDD1",
		000884 => x"E59F0340",
		000885 => x"EBFFFDCF",
		000886 => x"E59F033C",
		000887 => x"EBFFFDCD",
		000888 => x"E59F0338",
		000889 => x"EBFFFDCB",
		000890 => x"E59F0334",
		000891 => x"EBFFFDC9",
		000892 => x"E59F0330",
		000893 => x"EBFFFDC7",
		000894 => x"E59F032C",
		000895 => x"EBFFFDC5",
		000896 => x"E59F0328",
		000897 => x"EBFFFDC3",
		000898 => x"E59F0324",
		000899 => x"EBFFFDC1",
		000900 => x"E59F0320",
		000901 => x"EBFFFDBF",
		000902 => x"E59F031C",
		000903 => x"EBFFFDBD",
		000904 => x"E59F0318",
		000905 => x"EBFFFDBB",
		000906 => x"E59F0314",
		000907 => x"EBFFFDB9",
		000908 => x"E59F0310",
		000909 => x"EBFFFDB7",
		000910 => x"E59F030C",
		000911 => x"EBFFFDB5",
		000912 => x"E59F0308",
		000913 => x"EBFFFDB3",
		000914 => x"E59F0304",
		000915 => x"EBFFFDB1",
		000916 => x"E59F0300",
		000917 => x"EBFFFDAF",
		000918 => x"E59F02FC",
		000919 => x"EBFFFDAD",
		000920 => x"EAFFFEE0",
		000921 => x"E3A00069",
		000922 => x"EBFFFCD9",
		000923 => x"E59F02EC",
		000924 => x"EBFFFDA8",
		000925 => x"E59F02E8",
		000926 => x"EBFFFDA6",
		000927 => x"E59F02E4",
		000928 => x"EBFFFDA4",
		000929 => x"E59F02E0",
		000930 => x"EBFFFDA2",
		000931 => x"E59F02DC",
		000932 => x"EBFFFDA0",
		000933 => x"EAFFFED3",
		000934 => x"E20000FF",
		000935 => x"EBFFFCCC",
		000936 => x"E59F02CC",
		000937 => x"EBFFFD9B",
		000938 => x"EAFFFECE",
		000939 => x"E3A00072",
		000940 => x"EBFFFCC7",
		000941 => x"E3A006FF",
		000942 => x"E280F20F",
		000943 => x"EAFFFFFE",
		000944 => x"E3A00061",
		000945 => x"EBFFFCC2",
		000946 => x"E59F02A8",
		000947 => x"EBFFFD91",
		000948 => x"E59F02A4",
		000949 => x"EBFFFD8F",
		000950 => x"E59F02A0",
		000951 => x"EBFFFD8D",
		000952 => x"EAFFFEC0",
		000953 => x"E3A00066",
		000954 => x"EBFFFCB9",
		000955 => x"E59F0290",
		000956 => x"EBFFFD88",
		000957 => x"E59F028C",
		000958 => x"EBFFFD86",
		000959 => x"EAFFFEB9",
		000960 => x"E59F0284",
		000961 => x"EBFFFD83",
		000962 => x"E59F0280",
		000963 => x"EBFFFD81",
		000964 => x"EBFFFCA9",
		000965 => x"E3700001",
		000966 => x"0AFFFFFC",
		000967 => x"EBFFFCA6",
		000968 => x"E3700001",
		000969 => x"1AFFFFFC",
		000970 => x"E3A05000",
		000971 => x"E3A0C000",
		000972 => x"E1A02005",
		000973 => x"E1A01006",
		000974 => x"E3A03002",
		000975 => x"E3A00072",
		000976 => x"E58DC000",
		000977 => x"EBFFFCDE",
		000978 => x"E1A04000",
		000979 => x"EBFFFC9A",
		000980 => x"E3700001",
		000981 => x"E1A00004",
		000982 => x"1A00004E",
		000983 => x"E3540000",
		000984 => x"BAFFFFF1",
		000985 => x"EBFFFC9A",
		000986 => x"E3A03801",
		000987 => x"E2855001",
		000988 => x"E2433001",
		000989 => x"E1550003",
		000990 => x"1AFFFFEB",
		000991 => x"EAFFFEF4",
		000992 => x"E5DD1009",
		000993 => x"E3510042",
		000994 => x"1AFFFE92",
		000995 => x"E5DD000A",
		000996 => x"E3500052",
		000997 => x"1AFFFE8F",
		000998 => x"E3A04000",
		000999 => x"E5C43000",
		001000 => x"E1A00000",
		001001 => x"E5C42001",
		001002 => x"E1A00000",
		001003 => x"E5C41002",
		001004 => x"E1A00000",
		001005 => x"E5C40003",
		001006 => x"E1A00000",
		001007 => x"E241103E",
		001008 => x"E1A0000A",
		001009 => x"E1A02004",
		001010 => x"EBFFFD60",
		001011 => x"E5DD3007",
		001012 => x"E5C43004",
		001013 => x"E5DD2008",
		001014 => x"E5C42005",
		001015 => x"E5DD3009",
		001016 => x"E5C43006",
		001017 => x"E5DD200A",
		001018 => x"E1A0000A",
		001019 => x"E5C42007",
		001020 => x"EBFFFDAD",
		001021 => x"E3A03CFF",
		001022 => x"E28330FC",
		001023 => x"E1500003",
		001024 => x"E1A05000",
		001025 => x"8AFFFF48",
		001026 => x"E3700004",
		001027 => x"12844008",
		001028 => x"1280700B",
		001029 => x"0A000006",
		001030 => x"EBFFFC67",
		001031 => x"E3700001",
		001032 => x"0AFFFFFC",
		001033 => x"E1570004",
		001034 => x"E5C40000",
		001035 => x"E2844001",
		001036 => x"1AFFFFF8",
		001037 => x"E59F0158",
		001038 => x"EBFFFD36",
		001039 => x"E59F0154",
		001040 => x"EBFFFD34",
		001041 => x"E375000C",
		001042 => x"0A00000F",
		001043 => x"E3A04000",
		001044 => x"E285800C",
		001045 => x"E1A07004",
		001046 => x"E5D45000",
		001047 => x"E3A00077",
		001048 => x"E1A01006",
		001049 => x"E1A02007",
		001050 => x"E3A03002",
		001051 => x"E58D5000",
		001052 => x"EBFFFC93",
		001053 => x"E3500000",
		001054 => x"1AFFFFF7",
		001055 => x"E2844001",
		001056 => x"E1540008",
		001057 => x"E1A07004",
		001058 => x"1AFFFFF2",
		001059 => x"E59F0108",
		001060 => x"EBFFFD20",
		001061 => x"EAFFFE51",
		001062 => x"E59F0100",
		001063 => x"EBFFFD1D",
		001064 => x"EAFFFEAB",
		001065 => x"FFF011A4",
		001066 => x"FFF011F0",
		001067 => x"FFF01238",
		001068 => x"FFF01280",
		001069 => x"FFF012C8",
		001070 => x"FFF01310",
		001071 => x"FFF01358",
		001072 => x"FFF013C4",
		001073 => x"FFF013FC",
		001074 => x"FFF01460",
		001075 => x"FFF014C4",
		001076 => x"FFF0172C",
		001077 => x"FFF017D4",
		001078 => x"FFF01EE4",
		001079 => x"FFF01F14",
		001080 => x"FFF01514",
		001081 => x"FFF015AC",
		001082 => x"FFF015D4",
		001083 => x"FFF0161C",
		001084 => x"FFF01640",
		001085 => x"FFF016A4",
		001086 => x"FFF01690",
		001087 => x"FFF01588",
		001088 => x"FFF016D0",
		001089 => x"FFF0170C",
		001090 => x"FFF017F8",
		001091 => x"FFF01834",
		001092 => x"FFF019C0",
		001093 => x"FFF019DC",
		001094 => x"FFF019FC",
		001095 => x"FFF01A3C",
		001096 => x"FFF01A70",
		001097 => x"FFF01AAC",
		001098 => x"FFF01AE8",
		001099 => x"FFF01B0C",
		001100 => x"FFF01B48",
		001101 => x"FFF01B64",
		001102 => x"FFF01B7C",
		001103 => x"FFF01BC4",
		001104 => x"FFF01C04",
		001105 => x"FFF01C3C",
		001106 => x"FFF01C60",
		001107 => x"FFF01CA4",
		001108 => x"FFF01CE4",
		001109 => x"FFF01D10",
		001110 => x"FFF01D3C",
		001111 => x"FFF01D60",
		001112 => x"FFF01D88",
		001113 => x"FFF01DC0",
		001114 => x"FFF01DFC",
		001115 => x"FFF01E38",
		001116 => x"FFF01E78",
		001117 => x"FFF01EF0",
		001118 => x"FFF018DC",
		001119 => x"FFF01910",
		001120 => x"FFF0197C",
		001121 => x"FFF01E98",
		001122 => x"FFF01EC8",
		001123 => x"FFF01854",
		001124 => x"FFF01894",
		001125 => x"FFF0178C",
		001126 => x"FFF017A4",
		001127 => x"FFF017C4",
		001128 => x"FFF01F38",
		001129 => x"0D0A0D0A",
		001130 => x"0D0A2B2D",
		001131 => x"2D2D2D2D",
		001132 => x"2D2D2D2D",
		001133 => x"2D2D2D2D",
		001134 => x"2D2D2D2D",
		001135 => x"2D2D2D2D",
		001136 => x"2D2D2D2D",
		001137 => x"2D2D2D2D",
		001138 => x"2D2D2D2D",
		001139 => x"2D2D2D2D",
		001140 => x"2D2D2D2D",
		001141 => x"2D2D2D2D",
		001142 => x"2D2D2D2D",
		001143 => x"2D2D2D2D",
		001144 => x"2D2D2D2D",
		001145 => x"2D2D2D2D",
		001146 => x"2D2D2D2B",
		001147 => x"0D0A0000",
		001148 => x"7C202020",
		001149 => x"203C3C3C",
		001150 => x"2053544F",
		001151 => x"524D2043",
		001152 => x"6F726520",
		001153 => x"50726F63",
		001154 => x"6573736F",
		001155 => x"72205379",
		001156 => x"7374656D",
		001157 => x"202D2042",
		001158 => x"79205374",
		001159 => x"65706861",
		001160 => x"6E204E6F",
		001161 => x"6C74696E",
		001162 => x"67203E3E",
		001163 => x"3E202020",
		001164 => x"207C0D0A",
		001165 => x"00000000",
		001166 => x"2B2D2D2D",
		001167 => x"2D2D2D2D",
		001168 => x"2D2D2D2D",
		001169 => x"2D2D2D2D",
		001170 => x"2D2D2D2D",
		001171 => x"2D2D2D2D",
		001172 => x"2D2D2D2D",
		001173 => x"2D2D2D2D",
		001174 => x"2D2D2D2D",
		001175 => x"2D2D2D2D",
		001176 => x"2D2D2D2D",
		001177 => x"2D2D2D2D",
		001178 => x"2D2D2D2D",
		001179 => x"2D2D2D2D",
		001180 => x"2D2D2D2D",
		001181 => x"2D2D2D2D",
		001182 => x"2D2B0D0A",
		001183 => x"00000000",
		001184 => x"7C202020",
		001185 => x"20202020",
		001186 => x"20426F6F",
		001187 => x"746C6F61",
		001188 => x"64657220",
		001189 => x"666F7220",
		001190 => x"53544F52",
		001191 => x"4D20536F",
		001192 => x"43202020",
		001193 => x"56657273",
		001194 => x"696F6E3A",
		001195 => x"2031352E",
		001196 => x"30352E32",
		001197 => x"30313220",
		001198 => x"42202020",
		001199 => x"20202020",
		001200 => x"207C0D0A",
		001201 => x"00000000",
		001202 => x"7C202020",
		001203 => x"20202020",
		001204 => x"20202020",
		001205 => x"20202020",
		001206 => x"436F6E74",
		001207 => x"6163743A",
		001208 => x"2073746E",
		001209 => x"6F6C7469",
		001210 => x"6E674067",
		001211 => x"6F6F676C",
		001212 => x"656D6169",
		001213 => x"6C2E636F",
		001214 => x"6D202020",
		001215 => x"20202020",
		001216 => x"20202020",
		001217 => x"20202020",
		001218 => x"207C0D0A",
		001219 => x"00000000",
		001220 => x"2B2D2D2D",
		001221 => x"2D2D2D2D",
		001222 => x"2D2D2D2D",
		001223 => x"2D2D2D2D",
		001224 => x"2D2D2D2D",
		001225 => x"2D2D2D2D",
		001226 => x"2D2D2D2D",
		001227 => x"2D2D2D2D",
		001228 => x"2D2D2D2D",
		001229 => x"2D2D2D2D",
		001230 => x"2D2D2D2D",
		001231 => x"2D2D2D2D",
		001232 => x"2D2D2D2D",
		001233 => x"2D2D2D2D",
		001234 => x"2D2D2D2D",
		001235 => x"2D2D2D2D",
		001236 => x"2D2B0D0A",
		001237 => x"0D0A0000",
		001238 => x"203C2057",
		001239 => x"656C636F",
		001240 => x"6D652074",
		001241 => x"6F207468",
		001242 => x"65205354",
		001243 => x"4F524D20",
		001244 => x"536F4320",
		001245 => x"626F6F74",
		001246 => x"6C6F6164",
		001247 => x"65722063",
		001248 => x"6F6E736F",
		001249 => x"6C652120",
		001250 => x"3E0D0A20",
		001251 => x"3C205365",
		001252 => x"6C656374",
		001253 => x"20616E20",
		001254 => x"6F706572",
		001255 => x"6174696F",
		001256 => x"6E206672",
		001257 => x"6F6D2074",
		001258 => x"6865206D",
		001259 => x"656E7520",
		001260 => x"62656C6F",
		001261 => x"77206F72",
		001262 => x"20707265",
		001263 => x"7373203E",
		001264 => x"0D0A0000",
		001265 => x"203C2074",
		001266 => x"68652062",
		001267 => x"6F6F7420",
		001268 => x"6B657920",
		001269 => x"666F7220",
		001270 => x"696D6D65",
		001271 => x"64696174",
		001272 => x"65206170",
		001273 => x"706C6963",
		001274 => x"6174696F",
		001275 => x"6E207374",
		001276 => x"6172742E",
		001277 => x"203E0D0A",
		001278 => x"0D0A0000",
		001279 => x"2030202D",
		001280 => x"20626F6F",
		001281 => x"74206672",
		001282 => x"6F6D2063",
		001283 => x"6F726520",
		001284 => x"52414D20",
		001285 => x"28737461",
		001286 => x"72742061",
		001287 => x"70706C69",
		001288 => x"63617469",
		001289 => x"6F6E290D",
		001290 => x"0A203120",
		001291 => x"2D207072",
		001292 => x"6F677261",
		001293 => x"6D20636F",
		001294 => x"72652052",
		001295 => x"414D2076",
		001296 => x"69612055",
		001297 => x"4152545F",
		001298 => x"300D0A20",
		001299 => x"32202D20",
		001300 => x"636F7265",
		001301 => x"2052414D",
		001302 => x"2064756D",
		001303 => x"700D0A00",
		001304 => x"2033202D",
		001305 => x"20626F6F",
		001306 => x"74206672",
		001307 => x"6F6D2049",
		001308 => x"32432045",
		001309 => x"4550524F",
		001310 => x"4D0D0A20",
		001311 => x"34202D20",
		001312 => x"70726F67",
		001313 => x"72616D20",
		001314 => x"49324320",
		001315 => x"45455052",
		001316 => x"4F4D2076",
		001317 => x"69612055",
		001318 => x"4152545F",
		001319 => x"300D0A20",
		001320 => x"35202D20",
		001321 => x"73686F77",
		001322 => x"20636F6E",
		001323 => x"74656E74",
		001324 => x"206F6620",
		001325 => x"49324320",
		001326 => x"45455052",
		001327 => x"4F4D0D0A",
		001328 => x"00000000",
		001329 => x"2061202D",
		001330 => x"20617574",
		001331 => x"6F6D6174",
		001332 => x"69632062",
		001333 => x"6F6F7420",
		001334 => x"636F6E66",
		001335 => x"69677572",
		001336 => x"6174696F",
		001337 => x"6E0D0A20",
		001338 => x"68202D20",
		001339 => x"68656C70",
		001340 => x"0D0A2072",
		001341 => x"202D2072",
		001342 => x"65737461",
		001343 => x"72742073",
		001344 => x"79737465",
		001345 => x"6D0D0A0D",
		001346 => x"0A53656C",
		001347 => x"6563743A",
		001348 => x"20000000",
		001349 => x"0D0A0D0A",
		001350 => x"4170706C",
		001351 => x"69636174",
		001352 => x"696F6E20",
		001353 => x"77696C6C",
		001354 => x"20737461",
		001355 => x"72742061",
		001356 => x"75746F6D",
		001357 => x"61746963",
		001358 => x"616C6C79",
		001359 => x"20616674",
		001360 => x"65722064",
		001361 => x"6F776E6C",
		001362 => x"6F61642E",
		001363 => x"0D0A2D3E",
		001364 => x"20576169",
		001365 => x"74696E67",
		001366 => x"20666F72",
		001367 => x"20277374",
		001368 => x"6F726D5F",
		001369 => x"70726F67",
		001370 => x"72616D2E",
		001371 => x"62696E27",
		001372 => x"20696E20",
		001373 => x"62797465",
		001374 => x"2D737472",
		001375 => x"65616D20",
		001376 => x"6D6F6465",
		001377 => x"2E2E2E00",
		001378 => x"20455252",
		001379 => x"4F522120",
		001380 => x"50726F67",
		001381 => x"72616D20",
		001382 => x"66696C65",
		001383 => x"20746F6F",
		001384 => x"20626967",
		001385 => x"210D0A0D",
		001386 => x"0A000000",
		001387 => x"20496E76",
		001388 => x"616C6964",
		001389 => x"2070726F",
		001390 => x"6772616D",
		001391 => x"6D696E67",
		001392 => x"2066696C",
		001393 => x"65210D0A",
		001394 => x"0D0A5365",
		001395 => x"6C656374",
		001396 => x"3A200000",
		001397 => x"0D0A0D0A",
		001398 => x"41626F72",
		001399 => x"74206475",
		001400 => x"6D70696E",
		001401 => x"67206279",
		001402 => x"20707265",
		001403 => x"7373696E",
		001404 => x"6720616E",
		001405 => x"79206B65",
		001406 => x"792E0D0A",
		001407 => x"50726573",
		001408 => x"7320616E",
		001409 => x"79206B65",
		001410 => x"7920746F",
		001411 => x"20636F6E",
		001412 => x"74696E75",
		001413 => x"652E0D0A",
		001414 => x"0D0A0000",
		001415 => x"0D0A0D0A",
		001416 => x"44756D70",
		001417 => x"696E6720",
		001418 => x"636F6D70",
		001419 => x"6C657465",
		001420 => x"642E0D0A",
		001421 => x"0D0A5365",
		001422 => x"6C656374",
		001423 => x"3A200000",
		001424 => x"0D0A4170",
		001425 => x"706C6963",
		001426 => x"6174696F",
		001427 => x"6E207769",
		001428 => x"6C6C2073",
		001429 => x"74617274",
		001430 => x"20617574",
		001431 => x"6F6D6174",
		001432 => x"6963616C",
		001433 => x"6C792061",
		001434 => x"66746572",
		001435 => x"2075706C",
		001436 => x"6F61642E",
		001437 => x"0D0A2D3E",
		001438 => x"204C6F61",
		001439 => x"64696E67",
		001440 => x"20626F6F",
		001441 => x"7420696D",
		001442 => x"6167652E",
		001443 => x"2E2E0000",
		001444 => x"2055706C",
		001445 => x"6F616420",
		001446 => x"636F6D70",
		001447 => x"6C657465",
		001448 => x"0D0A0000",
		001449 => x"20496E76",
		001450 => x"616C6964",
		001451 => x"20626F6F",
		001452 => x"74206465",
		001453 => x"76696365",
		001454 => x"206F7220",
		001455 => x"66696C65",
		001456 => x"210D0A0D",
		001457 => x"0A53656C",
		001458 => x"6563743A",
		001459 => x"20000000",
		001460 => x"0D0A0D0A",
		001461 => x"456E7465",
		001462 => x"72206465",
		001463 => x"76696365",
		001464 => x"20616464",
		001465 => x"72657373",
		001466 => x"20283278",
		001467 => x"20686578",
		001468 => x"5F636861",
		001469 => x"72732C20",
		001470 => x"73657420",
		001471 => x"4C534220",
		001472 => x"746F2027",
		001473 => x"3027293A",
		001474 => x"20000000",
		001475 => x"0D0A496E",
		001476 => x"76616C69",
		001477 => x"64206164",
		001478 => x"64726573",
		001479 => x"73210D0A",
		001480 => x"0D0A5365",
		001481 => x"6C656374",
		001482 => x"3A200000",
		001483 => x"0D0A4461",
		001484 => x"74612077",
		001485 => x"696C6C20",
		001486 => x"6F766572",
		001487 => x"77726974",
		001488 => x"65205241",
		001489 => x"4D20636F",
		001490 => x"6E74656E",
		001491 => x"74210D0A",
		001492 => x"2D3E2057",
		001493 => x"61697469",
		001494 => x"6E672066",
		001495 => x"6F722027",
		001496 => x"73746F72",
		001497 => x"6D5F7072",
		001498 => x"6F677261",
		001499 => x"6D2E6269",
		001500 => x"6E272069",
		001501 => x"6E206279",
		001502 => x"74652D73",
		001503 => x"74726561",
		001504 => x"6D206D6F",
		001505 => x"64652E2E",
		001506 => x"2E000000",
		001507 => x"20446F77",
		001508 => x"6E6C6F61",
		001509 => x"6420636F",
		001510 => x"6D706C65",
		001511 => x"7465640D",
		001512 => x"0A000000",
		001513 => x"57726974",
		001514 => x"696E6720",
		001515 => x"62756666",
		001516 => x"65722074",
		001517 => x"6F206932",
		001518 => x"63204545",
		001519 => x"50524F4D",
		001520 => x"2E2E2E00",
		001521 => x"20436F6D",
		001522 => x"706C6574",
		001523 => x"65640D0A",
		001524 => x"0D0A0000",
		001525 => x"20496E76",
		001526 => x"616C6964",
		001527 => x"20626F6F",
		001528 => x"74206465",
		001529 => x"76696365",
		001530 => x"206F7220",
		001531 => x"66696C65",
		001532 => x"210D0A0D",
		001533 => x"0A000000",
		001534 => x"0D0A0D0A",
		001535 => x"456E7465",
		001536 => x"72206465",
		001537 => x"76696365",
		001538 => x"20616464",
		001539 => x"72657373",
		001540 => x"20283220",
		001541 => x"6865782D",
		001542 => x"63686172",
		001543 => x"732C2073",
		001544 => x"6574204C",
		001545 => x"53422074",
		001546 => x"6F202730",
		001547 => x"27293A20",
		001548 => x"00000000",
		001549 => x"20496E76",
		001550 => x"616C6964",
		001551 => x"20616464",
		001552 => x"72657373",
		001553 => x"210D0A0D",
		001554 => x"0A53656C",
		001555 => x"6563743A",
		001556 => x"20000000",
		001557 => x"0D0A0D0A",
		001558 => x"41626F72",
		001559 => x"74206475",
		001560 => x"6D70696E",
		001561 => x"67206279",
		001562 => x"20707265",
		001563 => x"7373696E",
		001564 => x"6720616E",
		001565 => x"79206B65",
		001566 => x"792E2049",
		001567 => x"66206E6F",
		001568 => x"20646174",
		001569 => x"61206973",
		001570 => x"2073686F",
		001571 => x"776E2C0D",
		001572 => x"0A000000",
		001573 => x"74686520",
		001574 => x"73656C65",
		001575 => x"63746564",
		001576 => x"20646576",
		001577 => x"69636520",
		001578 => x"6973206E",
		001579 => x"6F742072",
		001580 => x"6573706F",
		001581 => x"6E64696E",
		001582 => x"672E2050",
		001583 => x"72657373",
		001584 => x"20616E79",
		001585 => x"206B6579",
		001586 => x"20746F20",
		001587 => x"636F6E74",
		001588 => x"696E7565",
		001589 => x"2E0D0A0D",
		001590 => x"0A000000",
		001591 => x"0D0A0D0A",
		001592 => x"4175746F",
		001593 => x"6D617469",
		001594 => x"6320626F",
		001595 => x"6F742063",
		001596 => x"6F6E6669",
		001597 => x"67757261",
		001598 => x"74696F6E",
		001599 => x"20666F72",
		001600 => x"20706F77",
		001601 => x"65722D75",
		001602 => x"703A0D0A",
		001603 => x"00000000",
		001604 => x"5B333231",
		001605 => x"305D2063",
		001606 => x"6F6E6669",
		001607 => x"67757261",
		001608 => x"74696F6E",
		001609 => x"20444950",
		001610 => x"20737769",
		001611 => x"7463680D",
		001612 => x"0A203030",
		001613 => x"3030202D",
		001614 => x"20537461",
		001615 => x"72742062",
		001616 => x"6F6F746C",
		001617 => x"6F616465",
		001618 => x"7220636F",
		001619 => x"6E736F6C",
		001620 => x"650D0A20",
		001621 => x"30303031",
		001622 => x"202D2041",
		001623 => x"75746F6D",
		001624 => x"61746963",
		001625 => x"20626F6F",
		001626 => x"74206672",
		001627 => x"6F6D2063",
		001628 => x"6F726520",
		001629 => x"52414D0D",
		001630 => x"0A000000",
		001631 => x"20303031",
		001632 => x"30202D20",
		001633 => x"4175746F",
		001634 => x"6D617469",
		001635 => x"6320626F",
		001636 => x"6F742066",
		001637 => x"726F6D20",
		001638 => x"49324320",
		001639 => x"45455052",
		001640 => x"4F4D2028",
		001641 => x"41646472",
		001642 => x"65737320",
		001643 => x"30784130",
		001644 => x"290D0A0D",
		001645 => x"0A53656C",
		001646 => x"6563743A",
		001647 => x"20000000",
		001648 => x"0D0A0D0A",
		001649 => x"53544F52",
		001650 => x"4D20536F",
		001651 => x"4320626F",
		001652 => x"6F746C6F",
		001653 => x"61646572",
		001654 => x"0D0A0000",
		001655 => x"2730273A",
		001656 => x"20457865",
		001657 => x"63757465",
		001658 => x"2070726F",
		001659 => x"6772616D",
		001660 => x"20696E20",
		001661 => x"52414D2E",
		001662 => x"0D0A0000",
		001663 => x"2731273A",
		001664 => x"20577269",
		001665 => x"74652027",
		001666 => x"73746F72",
		001667 => x"6D5F7072",
		001668 => x"6F677261",
		001669 => x"6D2E6269",
		001670 => x"6E272074",
		001671 => x"6F207468",
		001672 => x"6520636F",
		001673 => x"72652773",
		001674 => x"2052414D",
		001675 => x"20766961",
		001676 => x"20554152",
		001677 => x"542E0D0A",
		001678 => x"00000000",
		001679 => x"2732273A",
		001680 => x"20507269",
		001681 => x"6E742063",
		001682 => x"75727265",
		001683 => x"6E742063",
		001684 => x"6F6E7465",
		001685 => x"6E74206F",
		001686 => x"6620636F",
		001687 => x"6D706C65",
		001688 => x"74652063",
		001689 => x"6F726520",
		001690 => x"52414D2E",
		001691 => x"0D0A0000",
		001692 => x"2733273A",
		001693 => x"204C6F61",
		001694 => x"6420626F",
		001695 => x"6F742069",
		001696 => x"6D616765",
		001697 => x"2066726F",
		001698 => x"6D204545",
		001699 => x"50524F4D",
		001700 => x"20616E64",
		001701 => x"20737461",
		001702 => x"72742061",
		001703 => x"70706C69",
		001704 => x"63617469",
		001705 => x"6F6E2E0D",
		001706 => x"0A000000",
		001707 => x"2734273A",
		001708 => x"20577269",
		001709 => x"74652027",
		001710 => x"73746F72",
		001711 => x"6D5F7072",
		001712 => x"6F677261",
		001713 => x"6D2E6269",
		001714 => x"6E272074",
		001715 => x"6F204932",
		001716 => x"43204545",
		001717 => x"50524F4D",
		001718 => x"20766961",
		001719 => x"20554152",
		001720 => x"542E0D0A",
		001721 => x"00000000",
		001722 => x"2735273A",
		001723 => x"20507269",
		001724 => x"6E742063",
		001725 => x"6F6E7465",
		001726 => x"6E74206F",
		001727 => x"66204932",
		001728 => x"43204545",
		001729 => x"50524F4D",
		001730 => x"2E0D0A00",
		001731 => x"2761273A",
		001732 => x"2053686F",
		001733 => x"77204449",
		001734 => x"50207377",
		001735 => x"69746368",
		001736 => x"20636F6E",
		001737 => x"66696775",
		001738 => x"72617469",
		001739 => x"6F6E7320",
		001740 => x"666F7220",
		001741 => x"6175746F",
		001742 => x"6D617469",
		001743 => x"6320626F",
		001744 => x"6F742E0D",
		001745 => x"0A000000",
		001746 => x"2768273A",
		001747 => x"2053686F",
		001748 => x"77207468",
		001749 => x"69732073",
		001750 => x"63726565",
		001751 => x"6E2E0D0A",
		001752 => x"00000000",
		001753 => x"2772273A",
		001754 => x"20526573",
		001755 => x"65742073",
		001756 => x"79737465",
		001757 => x"6D2E0D0A",
		001758 => x"0D0A0000",
		001759 => x"426F6F74",
		001760 => x"20454550",
		001761 => x"524F4D3A",
		001762 => x"20323478",
		001763 => x"786E6E6E",
		001764 => x"20286C69",
		001765 => x"6B652032",
		001766 => x"34414136",
		001767 => x"34292C20",
		001768 => x"37206269",
		001769 => x"74206164",
		001770 => x"64726573",
		001771 => x"73202B20",
		001772 => x"646F6E74",
		001773 => x"2D636172",
		001774 => x"65206269",
		001775 => x"742C0D0A",
		001776 => x"00000000",
		001777 => x"636F6E6E",
		001778 => x"65637465",
		001779 => x"6420746F",
		001780 => x"20493243",
		001781 => x"5F434F4E",
		001782 => x"54524F4C",
		001783 => x"4C45525F",
		001784 => x"302C206F",
		001785 => x"70657261",
		001786 => x"74696E67",
		001787 => x"20667265",
		001788 => x"7175656E",
		001789 => x"63792069",
		001790 => x"73203130",
		001791 => x"306B487A",
		001792 => x"2C0D0A00",
		001793 => x"6D617869",
		001794 => x"6D756D20",
		001795 => x"45455052",
		001796 => x"4F4D2073",
		001797 => x"697A6520",
		001798 => x"3D203635",
		001799 => x"35333620",
		001800 => x"62797465",
		001801 => x"203D3E20",
		001802 => x"31362062",
		001803 => x"69742061",
		001804 => x"64647265",
		001805 => x"73736573",
		001806 => x"2C0D0A00",
		001807 => x"66697865",
		001808 => x"6420626F",
		001809 => x"6F742064",
		001810 => x"65766963",
		001811 => x"65206164",
		001812 => x"64726573",
		001813 => x"733A2030",
		001814 => x"7841300D",
		001815 => x"0A0D0A00",
		001816 => x"5465726D",
		001817 => x"696E616C",
		001818 => x"20736574",
		001819 => x"75703A20",
		001820 => x"39363030",
		001821 => x"20626175",
		001822 => x"642C2038",
		001823 => x"20646174",
		001824 => x"61206269",
		001825 => x"74732C20",
		001826 => x"6E6F2070",
		001827 => x"61726974",
		001828 => x"792C2031",
		001829 => x"2073746F",
		001830 => x"70206269",
		001831 => x"740D0A0D",
		001832 => x"0A000000",
		001833 => x"466F7220",
		001834 => x"6D6F7265",
		001835 => x"20696E66",
		001836 => x"6F726D61",
		001837 => x"74696F6E",
		001838 => x"20736565",
		001839 => x"20746865",
		001840 => x"2053544F",
		001841 => x"524D2043",
		001842 => x"6F726520",
		001843 => x"2F205354",
		001844 => x"4F524D20",
		001845 => x"536F4320",
		001846 => x"64617461",
		001847 => x"73686565",
		001848 => x"740D0A00",
		001849 => x"68747470",
		001850 => x"3A2F2F6F",
		001851 => x"70656E63",
		001852 => x"6F726573",
		001853 => x"2E6F7267",
		001854 => x"2F70726F",
		001855 => x"6A656374",
		001856 => x"2C73746F",
		001857 => x"726D5F63",
		001858 => x"6F72650D",
		001859 => x"0A000000",
		001860 => x"68747470",
		001861 => x"3A2F2F6F",
		001862 => x"70656E63",
		001863 => x"6F726573",
		001864 => x"2E6F7267",
		001865 => x"2F70726F",
		001866 => x"6A656374",
		001867 => x"2C73746F",
		001868 => x"726D5F73",
		001869 => x"6F630D0A",
		001870 => x"00000000",
		001871 => x"436F6E74",
		001872 => x"6163743A",
		001873 => x"2073746E",
		001874 => x"6F6C7469",
		001875 => x"6E674067",
		001876 => x"6F6F676C",
		001877 => x"656D6169",
		001878 => x"6C2E636F",
		001879 => x"6D0D0A00",
		001880 => x"28632920",
		001881 => x"32303132",
		001882 => x"20627920",
		001883 => x"53746570",
		001884 => x"68616E20",
		001885 => x"4E6F6C74",
		001886 => x"696E670D",
		001887 => x"0A0D0A53",
		001888 => x"656C6563",
		001889 => x"743A2000",
		001890 => x"0D0A0D0A",
		001891 => x"496D6D65",
		001892 => x"72207765",
		001893 => x"6E6E2069",
		001894 => x"63682074",
		001895 => x"72617572",
		001896 => x"69672062",
		001897 => x"696E2C20",
		001898 => x"7472696E",
		001899 => x"6B206963",
		001900 => x"68206569",
		001901 => x"6E656E20",
		001902 => x"4B6F726E",
		001903 => x"2E0D0A00",
		001904 => x"57656E6E",
		001905 => x"20696368",
		001906 => x"2064616E",
		001907 => x"6E206E6F",
		001908 => x"63682074",
		001909 => x"72617572",
		001910 => x"69672062",
		001911 => x"696E2C20",
		001912 => x"7472696E",
		001913 => x"6B206963",
		001914 => x"68206E6F",
		001915 => x"63682765",
		001916 => x"6E204B6F",
		001917 => x"726E2E0D",
		001918 => x"0A000000",
		001919 => x"57656E6E",
		001920 => x"20696368",
		001921 => x"2044414E",
		001922 => x"4E206E6F",
		001923 => x"63682074",
		001924 => x"72617572",
		001925 => x"69672062",
		001926 => x"696E2C20",
		001927 => x"7472696E",
		001928 => x"6B206963",
		001929 => x"68204E4F",
		001930 => x"4348206E",
		001931 => x"656E204B",
		001932 => x"6F726E2E",
		001933 => x"0D0A0000",
		001934 => x"556E6420",
		001935 => x"77656E6E",
		001936 => x"20696368",
		001937 => x"2064616E",
		001938 => x"6E206E6F",
		001939 => x"63682074",
		001940 => x"72617572",
		001941 => x"69672062",
		001942 => x"696E2C20",
		001943 => x"66616E67",
		001944 => x"20696368",
		001945 => x"20616E20",
		001946 => x"766F6E20",
		001947 => x"766F726E",
		001948 => x"2E0D0A0D",
		001949 => x"0A000000",
		001950 => x"202D2048",
		001951 => x"65696E7A",
		001952 => x"20457268",
		001953 => x"61726474",
		001954 => x"0D0A0D0A",
		001955 => x"53656C65",
		001956 => x"63743A20",
		001957 => x"00000000",
		001958 => x"0D0A0D0A",
		001959 => x"5765276C",
		001960 => x"6C207365",
		001961 => x"6E642079",
		001962 => x"6F752062",
		001963 => x"61636B20",
		001964 => x"2D20746F",
		001965 => x"20746865",
		001966 => x"20667574",
		001967 => x"75726521",
		001968 => x"2E0D0A0D",
		001969 => x"0A000000",
		001970 => x"202D2044",
		001971 => x"6F63746F",
		001972 => x"7220456D",
		001973 => x"6D657420",
		001974 => x"4C2E2042",
		001975 => x"726F776E",
		001976 => x"0D0A0D0A",
		001977 => x"53656C65",
		001978 => x"63743A20",
		001979 => x"00000000",
		001980 => x"20496E76",
		001981 => x"616C6964",
		001982 => x"206F7065",
		001983 => x"72617469",
		001984 => x"6F6E210D",
		001985 => x"0A547279",
		001986 => x"20616761",
		001987 => x"696E3A20",
		001988 => x"00000000",
		001989 => x"0D0A0D0A",
		001990 => x"2D3E2053",
		001991 => x"74617274",
		001992 => x"696E6720",
		001993 => x"6170706C",
		001994 => x"69636174",
		001995 => x"696F6E2E",
		001996 => x"2E2E0D0A",
		001997 => x"0D0A0000",
		001998 => x"0D0A0D0A",
		001999 => x"41626F72",
		002000 => x"74656421",
		002001 => x"00000000",
		others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;